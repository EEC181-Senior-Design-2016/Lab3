module four_7hex (w,seg);

input [3:0] w;
output [0:6] seg;

assign seg[0] = (~w[3] & ~w[2] & ~w[1] & w[0]) |
	(~w[3] & w[2] & ~w[1] & ~w[0]) |
	(w[3] & ~w[2] & w[1] & w[0]) |
	(w[3] & w[2] & ~w[1] & w[0]);

assign seg[1] = (w[3] & w[1] & w[0]) |
	(w[2] & w[1] & ~w[0]) |
	(w[3] & w[2] & ~w[0]) |
	(~w[3] & w[2] & ~w[1] & w[0]);

assign seg[2] = (w[3] & w[2] & w[1]) |
	(w[3] & w[2] & ~w[0]) |
	(~w[3] & ~w[2] & w[1] & ~w[0]);

assign seg[3] = (w[2] & w[1] & w[0]) |
	(~w[3] & ~w[2] & ~w[1] & w[0]) |
	(~w[3] & w[2] & ~w[1] & ~w[0]) |
	(w[3] & ~w[2] & w[1] & ~w[0]);

assign seg[4] = (~w[3] & w[0]) |
	(~w[2] & ~w[1] & w[0]) |
	(~w[3] & w[2] & ~w[1]);

assign seg[5] = (~w[3] & w[1] & w[0]) |
	(~w[3] & ~w[2] & w[0]) |
	(~w[3] & ~w[2] & w[1]) |
	(w[3] & w[2] & ~w[1] & w[0]);

assign seg[6] = (~w[3] & ~w[2] & ~w[1]) |
	(~w[3] & w[2] & w[1] & w[0]) |
	(w[3] & w[2] & ~w[1] & ~w[0]);

endmodule